BZh91AY&SY_��� l_�Px����߰����P>r].��wFB�$�'�<A?T�Cj6���bdi��14��'�jhb=�F���4` H�M"Ci=L�z�zF�@ !�9�&& &#4���d�#RF��l������&�F �����?MȲVj�!a�?�A�`+���!|���)�6�%��8uG�� 7�jT�'<�p������2,_nb���LC��;cZ�*Ef<�0���8�[�,�3W{��$�� 9��w����}���)Lwm���
��t@v���a6�
�����;�,ڡ��Rh���k1�j4��h��S}�o�
I��S�(�2��4��+�$�l��ߑxp�6�{H��qZ�I���
[�Q��ezx�є]5#]#69"tAH��"�5GzWQ��D��W� {�g��/�	�؋+�=񛡼K,��r��Z�M���KT�
m�$�� j��g��ZL%����Oy�-��&g��,b3��K��UW� �������!�a��^�P�J�Yq=����J�y�7��]�c\�.�5%ႝ��Ɔ�%�E׎c(q5�o!�&20�E赨4q���K2�;`�rK	UV����EӅ3�����5�>\����%�Vp�u`��jr�z�^gpU�NW�R�����U��Ӥ�R�J�sC榿b�wl
�W}Hf�M}�#��K��gQ���D�ƛ�d�G��H��*�Y-9��/��d�����B~�w0U!���A���	��-"�sIl7	�Jo��K�hQ�&�Hv/�CL!��>"�"��Ȕ��&rZ�{mj���q��i�s��"�gtq����\�#�ۡ�:�]U1"Oi�Ө������W��A	���[AX�2�!�I��=%�����9�ؓ�	0xN�y�=���;=�ppl�0B�gJ���k0ц��Z�n��S33ad�M�3��V��hu@�L���\s�RMD̸:�'�l�}��Y��#���F��д~��H�
�x��